bhavana
sandrala
c
